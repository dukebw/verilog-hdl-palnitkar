module full_adder;
endmodule

module ripple_add;
    full_adder FullAdder0();
    full_adder FullAdder1();
    full_adder FullAdder2();
    full_adder FullAdder3();
endmodule
